-- stepmotor_tb.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity stepmotor_tb is
end entity stepmotor_tb;

architecture rtl of stepmotor_tb is
	component stepmotor is
		port (
			clk_clk            : in  std_logic                    := 'X'; -- clk
			leds_export        : out std_logic_vector(5 downto 0);        -- export
			reset_reset_n      : in  std_logic                    := 'X'; -- reset_n
			stepmotor_1_export : out std_logic_vector(3 downto 0)         -- export
		);
	end component stepmotor;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal stepmotor_inst_clk_bfm_clk_clk       : std_logic; -- stepmotor_inst_clk_bfm:clk -> [stepmotor_inst:clk_clk, stepmotor_inst_reset_bfm:clk]
	signal stepmotor_inst_reset_bfm_reset_reset : std_logic; -- stepmotor_inst_reset_bfm:reset -> stepmotor_inst:reset_reset_n

begin

	stepmotor_inst : component stepmotor
		port map (
			clk_clk            => stepmotor_inst_clk_bfm_clk_clk,       --         clk.clk
			leds_export        => open,                                 --        leds.export
			reset_reset_n      => stepmotor_inst_reset_bfm_reset_reset, --       reset.reset_n
			stepmotor_1_export => open                                  -- stepmotor_1.export
		);

	stepmotor_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => stepmotor_inst_clk_bfm_clk_clk  -- clk.clk
		);

	stepmotor_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => stepmotor_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => stepmotor_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of stepmotor_tb
